LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

BEGIN

Q <= Q + 1